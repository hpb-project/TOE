`timescale 1ns / 1ps
module bfifo #(
    	parameter RAM_STYLE  = "distributed",              // Specify RAM style: auto/block/distributed
	parameter DWID       = 18, 
	parameter AWID       = 6, 
	parameter AFULL_TH   = 4, 
	parameter AEMPTY_TH  = 4, 
	parameter DBG_WID    = 32 
) (
  //write clock domain
  input  		    clk,                          // write clock
  input 		    rst,                          // write reset
  input 		    wen,                           // Write enable
  input  [DWID-1:0]   	    wdata,                         // RAM input data
  output                    nfull,                         // 
  output                    nafull,                        // 
  output                    woverflow,                     // 
  output [AWID:0]           cnt_free,                      // the counter used in fifo for read clock domain 
  input                     ren,                           // Read Enable
  output [DWID-1:0]         rdata,                         // RAM output data
  output                    nempty,                        // 
  output                    naempty,                       // 
  output                    roverflow,                     // 
  output [AWID:0]           cnt_used ,                     // the counter used in fifo for write clock domain
  output [DBG_WID-1:0]      dbg_sig                        // debug signal
);


//////////////////////////////////////////////////////////////////////////////////
//  signal declare
//////////////////////////////////////////////////////////////////////////////////
wire                     old_ren        ;                     // Read Enable
wire  [DWID-1:0]         old_rdata      ;                     // RAM output data
wire                     old_nempty     ;                     // 
wire                     old_naempty    ;                     // 
wire                     old_roverflow  ;                     // 
 
//////////////////////////////////////////////////////////////////////////////////
//  old fifo
//////////////////////////////////////////////////////////////////////////////////
bfifo_reg #(
  .RAM_STYLE   ( RAM_STYLE   ),
  .DWID        ( DWID        ),
  .AWID        ( AWID        ),
  .AFULL_TH    ( AFULL_TH    ),
  .AEMPTY_TH   ( AEMPTY_TH   ),
  .DBG_WID     ( DBG_WID     )
) inst_fifo (
    .clk          ( clk          ),                 // write clock
    .rst          ( rst          ),                 // write reset
    .wen          ( wen           ),                 // Write enable
    .wdata        ( wdata         ),                 // RAM input data
    .nfull        ( nfull         ),                 // 
    .nafull       ( nafull        ),                 // 
    .woverflow    ( woverflow     ),                 // 
    .cnt_used     ( cnt_used      ),                 // the counter used in fifo for write clock domain
    .ren          ( old_ren       ),                 // Read Enable
    .rdata        ( old_rdata     ),                 // RAM output data
    .nempty       ( old_nempty    ),                 // 
    .naempty      ( naempty       ),                 // 
    .roverflow    ( old_roverflow ),                 // 
    .cnt_free     ( cnt_free      ),                 // the counter used in fifo for read clock domain 
    .dbg_sig      (               )                  // debug signal
);

//////////////////////////////////////////////////////////////////////////////////
//  new fifo read interface
//////////////////////////////////////////////////////////////////////////////////
fifo_rdif_tf #(
  .DWID        ( DWID ),
  .AWID        ( AWID )
) inst_fifo_rdif_tf (
  .clk               ( clk            ),                // Read clock
  .rst               ( rst            ),                // Read reset 
  .old_ren           ( old_ren        ),                // Read Enable
  .old_rdata         ( old_rdata      ),                // RAM output data
  .old_nempty        ( old_nempty     ),                // 
  .new_ren           ( ren            ),                // Read Enable
  .new_rdata         ( rdata          ),                // RAM output data
  .new_nempty        ( nempty         ),                // 
  .new_roverflow     ( roverflow      )                 // 
);

//////////////////////////////////////////////////////////////////////////////////
//  debug sig
//////////////////////////////////////////////////////////////////////////////////
assign dbg_sig = { 28'h0, woverflow, roverflow, nafull, nempty };

endmodule

module xilinx_simple_dual_port_2_clock_bram #(
  parameter RAM_WIDTH = 18,                       // Specify RAM data width
  parameter RAM_DEPTH = 1024,                     // Specify RAM depth (number of entires)
  //parameter RAM_PERFORMANCE = "HIGH_PERFORMANCE", // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
  parameter RAM_PERFORMANCE = "LOW_LATENCY", // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
  parameter INIT_FILE = ""                        // Specify name/location of RAM initialization file if using one (leave blank if not)
) (
  input [logb(RAM_DEPTH)-1:0] addra, // Write address bus, width determined from RAM_DEPTH
  input [logb(RAM_DEPTH)-1:0] addrb, // Read address bus, width determined from RAM_DEPTH
  input [RAM_WIDTH-1:0] dina,          // RAM input data
  input clka,                          // Write clock
  input clkb,                          // Read clock
  input wea,                           // Write enable
  input enb,                           // Read Enable, for additional power savings, disable when not in use
  input rstb,                          // Output reset (does not affect memory contents)
  input regceb,                        // Output register enable
  output [RAM_WIDTH-1:0] doutb         // RAM output data
);

  (* ram_extract="yes", ram_style="block" *) reg [RAM_WIDTH-1:0] BRAM [RAM_DEPTH-1:0];
  reg [RAM_WIDTH-1:0] ram_data = {RAM_WIDTH{1'b0}};

  // The folowing code either initializes the memory values to a specified file or to all zeros to match hardware
  generate
    if (INIT_FILE != "") begin: use_init_file
      initial
        $readmemh(INIT_FILE, BRAM, 0, RAM_DEPTH-1);
    end else begin: init_bram_to_zero
      integer ram_index;
      initial
        for (ram_index = 0; ram_index < RAM_DEPTH; ram_index = ram_index + 1)
          BRAM[ram_index] = {RAM_WIDTH{1'b0}};
    end
  endgenerate

  always @(posedge clka)
    if (wea)
      BRAM[addra] <= dina; 
       
  always @(posedge clkb)
    if (enb)
      ram_data <= BRAM[addrb];

  //  The following code generates HIGH_PERFORMANCE (use output register) or LOW_LATENCY (no output register)
  generate
    if (RAM_PERFORMANCE == "LOW_LATENCY") begin: no_output_register

      // The following is a 1 clock cycle read latency at the cost of a longer clock-to-out timing
       assign doutb = ram_data;

    end else begin: output_register

      // The following is a 2 clock cycle read latency with improve clock-to-out timing

      reg [RAM_WIDTH-1:0] doutb_reg = {RAM_WIDTH{1'b0}};

      always @(posedge clkb)
        if (rstb)
          doutb_reg <= {RAM_WIDTH{1'b0}};
        else if (regceb)
          doutb_reg <= ram_data;

      assign doutb = doutb_reg;

    end
  endgenerate

//  The following function calculates the address width based on specified RAM depth
function integer logb;
  input integer depth;
  integer depth_reg;
	begin
        depth_reg = depth;
        for (logb=0; depth_reg>0; logb=logb+1)begin
          depth_reg = depth_reg >> 1;
        end
        if( 2**logb >= depth*2 )begin
          logb = logb - 1;
        end
	end 
endfunction

endmodule

//  Xilinx Simple Dual Port Single Clock RAM
//  This code implements a paramtizable SDP single clock memory.
//  If a reset or enable is not necessary, it may be tied off or removed from the code.

module xilinx_simple_dual_port_1_clock_bram #(
  parameter RAM_WIDTH = 18,                       // Specify RAM data width
  parameter RAM_DEPTH = 1024,                     // Specify RAM depth (number of entires)
  //parameter RAM_PERFORMANCE = "HIGH_PERFORMANCE", // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
  parameter RAM_PERFORMANCE = "LOW_LATENCY", // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
  parameter INIT_FILE = ""                        // Specify name/location of RAM initialization file if using one (leave blank if not)
) (
  input [logb(RAM_DEPTH)-1:0] addra, // Write address bus, width determined from RAM_DEPTH
  input [logb(RAM_DEPTH)-1:0] addrb, // Read address bus, width determined from RAM_DEPTH
  input [RAM_WIDTH-1:0] dina,          // RAM input data
  input clka,                          // Clock
  input wea,                           // Write enable
  input enb,                           // Read Enable, for additional power savings, disable when not in use
  input rstb,                          // Output reset (does not affect memory contents)
  input regceb,                        // Output register enable
  output [RAM_WIDTH-1:0] doutb         // RAM output data
);

  (* ram_extract="yes", ram_style="block" *) reg [RAM_WIDTH-1:0] BRAM [RAM_DEPTH-1:0];
  reg [RAM_WIDTH-1:0] ram_data = {RAM_WIDTH{1'b0}};

  // The folowing code either initializes the memory values to a specified file or to all zeros to match hardware
  generate
    if (INIT_FILE != "") begin: use_init_file
      initial begin
        $readmemh(INIT_FILE, BRAM, 0, RAM_DEPTH-1);
      end
	/* synthesis translate_off */ 
      initial begin
	$display("INIT_FILE=%s", INIT_FILE);
      end
	/* synthesis translate_on */ 
    end else begin: init_bram_to_zero
      integer ram_index;
      initial
        for (ram_index = 0; ram_index < RAM_DEPTH; ram_index = ram_index + 1)
          BRAM[ram_index] = {RAM_WIDTH{1'b0}};
    end
  endgenerate

  always @(posedge clka) begin
    if (wea)
      BRAM[addra] <= dina; 
    if (enb)
      ram_data <= BRAM[addrb];
  end        

  //  The following code generates HIGH_PERFORMANCE (use output register) or LOW_LATENCY (no output register)
  generate
    if (RAM_PERFORMANCE == "LOW_LATENCY") begin: no_output_register

      // The following is a 1 clock cycle read latency at the cost of a longer clock-to-out timing
       assign doutb = ram_data;

    end else begin: output_register

      // The following is a 2 clock cycle read latency with improve clock-to-out timing

      reg [RAM_WIDTH-1:0] doutb_reg = {RAM_WIDTH{1'b0}};

      always @(posedge clka)
        if (rstb)
          doutb_reg <= {RAM_WIDTH{1'b0}};
        else if (regceb)
          doutb_reg <= ram_data;

      assign doutb = doutb_reg;

    end
  endgenerate

//  The following function calculates the address width based on specified RAM depth
function integer logb;
  input integer depth;
  integer depth_reg;
	begin
        depth_reg = depth;
        for (logb=0; depth_reg>0; logb=logb+1)begin
          depth_reg = depth_reg >> 1;
        end
        if( 2**logb >= depth*2 )begin
          logb = logb - 1;
        end
	end 
endfunction

endmodule


//  Xilinx Simple Dual Port 2 Clock RAM
//  This code implements a paramtizable SDP dual clock memory.
//  If a reset or enable is not necessary, it may be tied off or removed from the code.

module xilinx_simple_dual_port_2_clock_dram #(
  parameter RAM_WIDTH = 18,                       // Specify RAM data width
  parameter RAM_DEPTH = 1024,                     // Specify RAM depth (number of entires)
  //parameter RAM_PERFORMANCE = "HIGH_PERFORMANCE", // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
  parameter RAM_PERFORMANCE = "LOW_LATENCY", // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
  parameter INIT_FILE = ""                        // Specify name/location of RAM initialization file if using one (leave blank if not)
) (
  input [logb(RAM_DEPTH)-1:0] addra, // Write address bus, width determined from RAM_DEPTH
  input [logb(RAM_DEPTH)-1:0] addrb, // Read address bus, width determined from RAM_DEPTH
  input [RAM_WIDTH-1:0] dina,          // RAM input data
  input clka,                          // Write clock
  input clkb,                          // Read clock
  input wea,                           // Write enable
  input enb,                           // Read Enable, for additional power savings, disable when not in use
  input rstb,                          // Output reset (does not affect memory contents)
  input regceb,                        // Output register enable
  output [RAM_WIDTH-1:0] doutb         // RAM output data
);

  (* ram_extract="yes", ram_style="distributed" *) reg [RAM_WIDTH-1:0] BRAM [RAM_DEPTH-1:0];
  reg [RAM_WIDTH-1:0] ram_data = {RAM_WIDTH{1'b0}};

  // The folowing code either initializes the memory values to a specified file or to all zeros to match hardware
  generate
    if (INIT_FILE != "") begin: use_init_file
      initial
        $readmemh(INIT_FILE, BRAM, 0, RAM_DEPTH-1);
    end else begin: init_bram_to_zero
      integer ram_index;
      initial
        for (ram_index = 0; ram_index < RAM_DEPTH; ram_index = ram_index + 1)
          BRAM[ram_index] = {RAM_WIDTH{1'b0}};
    end
  endgenerate

  always @(posedge clka)
    if (wea)
      BRAM[addra] <= dina; 
       
  always @(posedge clkb)
    if (enb)
      ram_data <= BRAM[addrb];

  //  The following code generates HIGH_PERFORMANCE (use output register) or LOW_LATENCY (no output register)
  generate
    if (RAM_PERFORMANCE == "LOW_LATENCY") begin: no_output_register

      // The following is a 1 clock cycle read latency at the cost of a longer clock-to-out timing
       assign doutb = ram_data;

    end else begin: output_register

      // The following is a 2 clock cycle read latency with improve clock-to-out timing

      reg [RAM_WIDTH-1:0] doutb_reg = {RAM_WIDTH{1'b0}};

      always @(posedge clkb)
        if (rstb)
          doutb_reg <= {RAM_WIDTH{1'b0}};
        else if (regceb)
          doutb_reg <= ram_data;

      assign doutb = doutb_reg;

    end
  endgenerate

//  The following function calculates the address width based on specified RAM depth
function integer logb;
  input integer depth;
  integer depth_reg;
	begin
        depth_reg = depth;
        for (logb=0; depth_reg>0; logb=logb+1)begin
          depth_reg = depth_reg >> 1;
        end
        if( 2**logb >= depth*2 )begin
          logb = logb - 1;
        end
	end 
endfunction

endmodule